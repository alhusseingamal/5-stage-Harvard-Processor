LIBRARY IEEE;
USE IEEE.STD_LOGIC_1164.ALL;
USE IEEE.numeric_std.all;

entity ID_EX_reg is
    port (
        clk : in std_logic;
        reset, flush : in std_logic;
        WB_in : IN std_logic_vector(1 downto 0);
        WB_out : OUT std_logic_vector(1 downto 0);
        RegRead_in : IN std_logic_vector(1 downto 0);
        RegRead_out : OUT std_logic_vector(1 downto 0);
        is_imm_in: IN std_logic;
        is_imm_out: OUT std_logic;
        MemtoReg_in : IN std_logic;
        MemtoReg_out : OUT std_logic;
        MemWrite_in : IN std_logic;
        MemWrite_out : OUT std_logic;
        MemRead_in : IN std_logic;
        MemRead_out : OUT std_logic;
        AluSrc_in : IN std_logic;
        AluSrc_out : OUT std_logic;
        ALUOp_in : IN std_logic_vector(3 downto 0);
        ALUOp_out : OUT std_logic_vector(3 downto 0);
        Predicted_in : IN std_logic;
        Predicted_out : OUT std_logic;
        branch_in : IN std_logic;
        branch_out : OUT std_logic;
        jmp_in : IN std_logic;
        jmp_out : OUT std_logic;
        Protect_in : IN std_logic;
        Protect_out : OUT std_logic;
        Free_in : IN std_logic;
        Free_out : OUT std_logic;
        i_RET : IN std_logic;
        o_RET : OUT std_logic;
        i_RTI : IN std_logic;
        o_RTI : OUT std_logic;
        i_popCCR : IN std_logic;
        o_popCCR : OUT std_logic;
        stack_op_in : IN std_logic;
        stack_op_out : OUT std_logic;
        push_pop_in : IN std_logic;
        push_pop_out : OUT std_logic;
        PC_data_mem_sel_in : IN std_logic;
        PC_data_mem_sel_out : OUT std_logic;
        Rsrc2_data_mem_sel_in : IN std_logic;
        Rsrc2_data_mem_sel_out : OUT std_logic;
        CCR_data_mem_sel_in : IN std_logic;
        CCR_data_mem_sel_out : OUT std_logic;
        STD_data_mem_sel_in : IN std_logic;
        STD_data_mem_sel_out : OUT std_logic;
        swap_in : IN std_logic;
        swap_out : OUT std_logic;
        src1_in : IN std_logic_vector(31 downto 0);
        src1_out : OUT std_logic_vector(31 downto 0);
        src2_in : IN std_logic_vector(31 downto 0);
        src2_out : OUT std_logic_vector(31 downto 0);
        STD_in : IN std_logic_vector(31 downto 0);
        STD_out : OUT std_logic_vector(31 downto 0);
        PC_in : IN std_logic_vector(31 downto 0);
        PC_out : OUT std_logic_vector(31 downto 0);
        Rs_in : IN std_logic_vector(2 downto 0);
        Rs_out : OUT std_logic_vector(2 downto 0);
        Rt_in : IN std_logic_vector(2 downto 0);
        Rt_out : OUT std_logic_vector(2 downto 0);
        Rd_in : IN std_logic_vector(2 downto 0);
        Rd_out : OUT std_logic_vector(2 downto 0);
        OutPortSignal_in : IN std_logic;
        OutPortSignal_out : OUT std_logic 
    );
end ID_EX_reg;

architecture Behavioral of ID_EX_reg is

begin
    process(clk, reset)
    begin
        if reset = '1' then
            WB_out <= (others => '0');
            RegRead_out <= (others => '0');
            is_imm_out <= '0';
            MemtoReg_out <= '0';
            MemWrite_out <= '0';
            MemRead_out <= '0';
            AluSrc_out <= '0';
            ALUOp_out <= (others => '1');
            Predicted_out <= '0';
            branch_out <= '0';
            jmp_out <= '0';
            o_RET <= '0';
            o_RTI <= '0';
            o_popCCR <= '0';
            stack_op_out <= '0';
            push_pop_out <= '0';
            PC_data_mem_sel_out <= '0';
            Rsrc2_data_mem_sel_out <= '0';
            CCR_data_mem_sel_out <= '0';
            STD_data_mem_sel_out <= '0';
            swap_out <= '0';
            src1_out <= (others => '0');
            src2_out <= (others => '0');
            STD_out <= (others => '0');
            PC_out <= (others => '0');
            Rs_out <= (others => '0');
            Rt_out <= (others => '0');
            Rd_out <= (others => '0');
            OutPortSignal_out <= '0';
            Protect_out <= '0';
            Free_out <= '0';
        elsif falling_edge(clk) then
            if flush = '1' then
                WB_out <= (others => '0');
                RegRead_out <= (others => '0');
                is_imm_out <= '0';
                MemtoReg_out <= '0'; 
                MemWrite_out <= '0';
                MemRead_out <= '0';
                AluSrc_out <= '0';
                ALUOp_out <= (others => '1');
                Predicted_out <= '0';
                branch_out <= '0';
                jmp_out <= '0';
                o_RET <= '0';
                o_RTI <= '0';
                o_popCCR <= '0';
                stack_op_out <= '0';
                push_pop_out <= '0';
                PC_data_mem_sel_out <= '0';
                Rsrc2_data_mem_sel_out <= '0';
                CCR_data_mem_sel_out <= '0';
                STD_data_mem_sel_out <= '0';
                swap_out <= '0';
                src1_out <= (others => '0');
                src2_out <= (others => '0');
                STD_out <= (others => '0');
                PC_out <= (others => '0');
                Rs_out <= (others => '0');
                Rt_out <= (others => '0');
                Rd_out <= (others => '0');
                OutPortSignal_out <= '0';
                Protect_out <= '0';
                Free_out <= '0';
            else
                is_imm_out <= is_imm_in;
                WB_out <= WB_in;
                RegRead_out <= RegRead_in;
                MemtoReg_out <= MemtoReg_in;
                MemWrite_out <= MemWrite_in;
                MemRead_out <= MemRead_in;
                AluSrc_out <= AluSrc_in;
                ALUOp_out <= ALUOp_in;
                Predicted_out <= Predicted_in;
                branch_out <= branch_in;
                jmp_out <= jmp_in;
                Protect_out <= Protect_in;
                Free_out <= Free_in;
                o_RET <= i_RET;
                o_RTI <= i_RTI;
                o_popCCR <= i_popCCR;
                stack_op_out <= stack_op_in;
                push_pop_out <= push_pop_in;
                PC_data_mem_sel_out <= PC_data_mem_sel_in;
                Rsrc2_data_mem_sel_out <= Rsrc2_data_mem_sel_in;
                CCR_data_mem_sel_out <= CCR_data_mem_sel_in;
                STD_data_mem_sel_out <= STD_data_mem_sel_in;
                swap_out <= swap_in;
                src1_out <= src1_in;
                src2_out <= src2_in;
                STD_out <= STD_in;
                PC_out <= PC_in;
                Rs_out <= Rs_in;
                Rt_out <= Rt_in;
                Rd_out <= Rd_in;
                OutPortSignal_out <= OutPortSignal_in;
            end if;
        end if;
    end process;

end Behavioral;